module top(
    input [15:0] sw,
    input btnC, // Clock
    input btnU, // Reset
    output [15:0] led, // A & B display
    output [6:0] seg,
    output [3:0] an
);

endmodule
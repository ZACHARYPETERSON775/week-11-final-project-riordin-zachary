module memory(
    input [7:0] data,
    input store,
    output reg [7:0] mem
);

    
endmodule